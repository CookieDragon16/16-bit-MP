library verilog;
use verilog.vl_types.all;
entity ERM16_tb is
end ERM16_tb;
