library verilog;
use verilog.vl_types.all;
entity tb_alu16 is
end tb_alu16;
